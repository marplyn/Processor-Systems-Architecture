module rom256_32 (          // создать блок с именем rom256_32
  input   [31:0]   A,     // 32-битный адресный вход
  
  output  [31:0]   RD     // 32-битный выход считанных данных
);

    reg [31:0] RAM [0:255];   // создать память с 256-ю 32-битными ячейками

    initial $readmemh("mem.txt", RAM);  // поместить при запуске микросхемы в
                                      // память RAM содержимое файла mem.txt


    assign RD = RAM[A];   // реализация порта на чтение


endmodule                 //  конец описания модуля