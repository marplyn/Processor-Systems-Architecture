module tb_rom;

reg   [31:0] adr;                      // создаем регистр для управления входом адреса
wire  [255:0] rd;                       // создаем провод для подключения к выходу памяти

rom256_32 dut (.A(adr), .RD(rd));        // подключаем проверяемый модуль

integer         i;                      // переменная для цикла for
integer         file_mem;               // для сохранения дескриптора файла
reg     [255:0] new_data;               // для сохранения очередного значения из файла

initial
  file_mem = $fopen("mem.txt", "r");  // получение дескриптора файла для последующего чтения "r"

initial begin
  for (i = 0; i < 31; i = i + 1) begin // подобно синтаксису C - выполнить цикл 8 раз для i от 0 до 7
    adr = i;                          // подать на вход адреса текущее значение i
    $fscanf(file_mem, "%b", new_data);// считать очередную строку (одно значение) из файла в new_data 
    #10;                              // задержка 10 единиц времени симуляции
    if (new_data != rd) begin         // если значение выдаваемое блоком памяти не равно значению из файла, то
      $display($time, "BAD!  adr = %d, file = %h, memory = %h", adr, new_data, rd);  // сообщить об ошибке
    end                              
  end
  $fclose(file_mem);                  // закрыть файл
  $finish;                            // закончить симуляцию
end

endmodule